// Defines for EDU-FPGA
`define PMOD0
`define PMOD1
`define ARDUINO
