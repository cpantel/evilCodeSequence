// Defines for EDU-FPGA
`define noPMOD0_DEV
`define noPMOD1_DEV
`define ARDUINO_DEV
`define RTC_DEV
`define noSERVO_DEV
`define UART_DEV

`define noPMOD0_CONN
`define noPMOD1_CONN
`define ARDUINO_CONN

