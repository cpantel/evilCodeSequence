// Defines for EDU-FPGA
`define noPMOD0_DEV
`define noPMOD1_DEV
`define noARDUINO_DEV

`define noPMOD0_CONN
`define noPMOD1_CONN
`define ARDUINO_CONN
