// Defines for servo_device running in EDU-FPGA
`define RTC_DEV
`define SERVO_DEV
`define UART_DEV

`define ARDUINO_CONN

