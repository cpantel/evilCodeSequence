// Defines for EDU-FPGA
`define noPMOD0_DEV
`define noPMOD1_DEV
`define noARDUINO_DEV
`define RTC_DEV
`define noSERVO_DEV
`define UART_DEV
`define KITT_DEV
`define noSEQUENCER_DEV

`define PMOD0_CONN
`define noPMOD1_CONN
`define noARDUINO_CONN

