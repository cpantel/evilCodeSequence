// Defines for EDU-FPGA
`define noPMOD0_DEV
`define noPMOD1_DEV
`define noARDUINO_DEV
`define RTC_DEV
`define SERVO_DEV
`define UART_DEV
`define PWM_DEV

`define KITT_DEV
`define SEQUENCER_DEV

`define PMOD0_CONN
`define noPMOD1_CONN
`define ARDUINO_CONN

