// Defines for EDU-FPGA
`define PMOD0_DEV
`define PMOD1_DEV
`define ARDUINO_DEV
`define noRTC_DEV
`define noSERVO_DEV
`define UART_DEV

`define PMOD0_CONN
`define PMOD1_CONN
`define ARDUINO_CONN

