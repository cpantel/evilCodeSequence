// Defines for EDU-FPGA
`define PMOD0_DEV
`define noPMOD1_DEV
`define noARDUINO_DEV
`define noRTC_DEV
`define noSERVO_DEV
`define UART_DEV

`define PMOD0_CONN
`define noPMOD1_CONN
`define noARDUINO_CONN

