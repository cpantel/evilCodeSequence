// Defines for servo_device running in EDU-FPGA
`define noPMOD0_DEV
`define noPMOD1_DEV
`define noARDUINO_DEV
`define noRTC_DEV
`define SERVO_DEV
`define UART_DEV

`define noPMOD0_CONN
`define noPMOD1_CONN
`define ARDUINO_CONN

