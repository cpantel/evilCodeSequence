// Defines for EDU-FPGA
`define noPMOD0
`define noPMOD1
`define noARDUINO
