// Defines for EDU-FPGA
`define noPMOD0_DEV
`define noPMOD1_DEV
`define noARDUINO_DEV
`define RTC_DEV
`define noSERVO_DEV
`define UART_DEV
`define noKITT_DEV
`define noSEQUENCER_DEV

`define noPMOD0_CONN
`define noPMOD1_CONN
`define noARDUINO_CONN

