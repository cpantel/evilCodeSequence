// Defines for kitt running in EDU-FPGA
`define KITT_DEV
`define UART_DEV

`define PMOD0_CONN


