// Valid defines for EDU-FPGA
//
// `define PMOD0_DEV
// `define PMOD1_DEV
// `define ARDUINO_DEV
// `define RTC_DEV
// `define SERVO_DEV
// `define KITT_DEV
// `define UART_DEV
//
// `define PMOD0_CONN
// `define PMOD1_CONN
// `define ARDUINO_CONN

